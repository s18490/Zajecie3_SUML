��X(      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.0.1�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�auto�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�objawy��wiek��choroby��wzrost�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��h2�f8�����R�(KhHNNNJ����J����K t�b�C              �?�t�bhLh&�scalar���hGC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hK�
node_count�K�nodes�h(h+K ��h-��R�(KK��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hxhGK ��hyhGK��hzhGK��h{hXK��h|hXK ��h}hGK(��h~hXK0��uK8KKt�b�B                              @��W3�?,            �Q@                           @��<D�m�?            �H@������������������������       �                     G@������������������������       �                     @������������������������       �                     6@�t�b�values�h(h+K ��h-��R�(KKKK��hX�CP      G@      9@      G@      @      G@                      @              6@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                              @:%�[��?,            �Q@                            @8��8���?             H@������������������������       �                     B@                          �g@�q�q�?             (@                          �@@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     7@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�     �E@      <@     �E@      @      B@              @      @      �?      @      �?                      @      @                      7@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @.}Z*�?)            �Q@                            @�nkK�?             G@������������������������       �                    �C@                          Pf@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     9@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      F@      ;@      F@       @     �C@              @       @               @      @                      9@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�C�                            @`��_��?,            �Q@������������������������       �                     B@������������������������       �                    �A@�t�bh�h(h+K ��h-��R�(KKKK��hX�C0      B@     �A@      B@                     �A@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoK	hph(h+K ��h-��R�(KK	��hw�B�                              @L�];�?+            �Q@������������������������       �                    �A@                            @r�q��?             B@                        0E�G@      �?             (@                          �g@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     8@�t�bh�h(h+K ��h-��R�(KK	KK��hX�C�     �D@      >@     �A@              @      >@      @      @      @       @               @      @                      @              8@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�Bh                            �d@.}Z*�?+            �Q@                           @�IєX�?
             1@������������������������       �        	             0@������������������������       �                     �?                            @|��?���?!             K@������������������������       �                     ;@       
                   �0@ 7���B�?             ;@       	                     @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     7@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      F@      ;@      0@      �?      0@                      �?      <@      :@      ;@              �?      :@      �?      @      �?                      @              7@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                            �E@�J�T�?(            �Q@                            @���V��?            �F@������������������������       �                     C@������������������������       �                     @                            @�n_Y�K�?             :@������������������������       �                     $@������������������������       �                     0@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp      H@      7@      C@      @      C@                      @      $@      0@      $@                      0@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @R_u^|�?/            �Q@                           @�C��2(�?             F@                            @Du9iH��?            �E@������������������������       �                    �@@       
                   �g@�z�G��?             $@                           �?      �?             @������������������������       �                      @       	                   �@@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     ;@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      D@      ?@      D@      @      D@      @     �@@              @      @      @      @       @              �?      @      �?                      @      @                      �?              ;@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ	�tlhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                            �d@DX�\��?.            �Q@                            @@4և���?             ,@������������������������       �        
             *@������������������������       �                     �?                            @6C�z��?#            �L@������������������������       �                     8@                            @6YE�t�?            �@@       	                   �@@�q�q�?             (@������������������������       �                     @
                          �g@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     5@�t�bh�h(h+K ��h-��R�(KKKK��hX�C�      E@      =@      *@      �?      *@                      �?      =@      <@      8@              @      <@      @      @      @               @      @              @       @                      5@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ޡhG        hNhG        h>Kh?Kh@h(h+K ��h-��R�(KK��hX�C              �?�t�bhLh]hGC       ���R�haKhbheKh(h+K ��h-��R�(KK��hG�C       �t�bK��R�}�(hKhoKhph(h+K ��h-��R�(KK��hw�B�                              @"` Y��?*            �Q@������������������������       �                    �D@                          @@@�r����?             >@                            @���|���?             &@������������������������       �                     @������������������������       �                     @������������������������       �                     3@�t�bh�h(h+K ��h-��R�(KKKK��hX�Cp     �F@      :@     �D@              @      :@      @      @      @                      @              3@�t�bubhhubehhub.